module friscv_uc(
    
);
endmodule