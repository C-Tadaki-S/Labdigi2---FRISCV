module friscv(

    // Entradas
    input               clock,              // Clock do circuito
    input               reset,              // Reseta o circuito
    input               liga_suco_1,        // Entrada do botão que ativa para o suco 1
    input               liga_suco_1,        // Entrada do botão que ativa para o suco 2

    // Saídas

    // Saídas de depuração
);



endmodule